library verilog;
use verilog.vl_types.all;
entity MIPSdatapath_testbench is
end MIPSdatapath_testbench;
